///////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////sequencer///////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//import UART_Package::*;
/*
class My_Sequencer extends uvm_sequencer #(Radwa_sequence_item);

      `uvm_component_utils (My_Sequencer)
///////////////////////////////////////////////new/////////////////////////////////////////////////////////////
  function new (string name, uvm_component parent);
     super.new(name, parent);
  endfunction


//////////////////////////////////////////build_phase//////////////////////////////////////////////////////////
    function void build_phase(uvm_phase phase);
       super.build_phase(phase);
       $display("build phase of sequencer");
    endfunction


///////////////////////////////////////////connect_phase///////////////////////////////////////////////////////
    function void connect_phase(uvm_phase phase);
       super.connect_phase(phase);
       $display("connect phase of sequencer");
    endfunction


//////////////////////////////////////////////run_phase////////////////////////////////////////////////////////
    task run_phase(uvm_phase phase);
       super.run_phase(phase);
       $display("run phase of sequencer");
    endtask
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
endclass
*/