///////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////Agent///////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////

class Agent_IN extends uvm_agent;

  `uvm_component_utils (Agent_IN)
  
  Radwa_monitor_in Rad_mon_in;
  ///////////tlm
  uvm_analysis_port #(Radwa_sequence_item) My_analysis_port;
  
  virtual INTF_UART U_intf;
///////////////////////////////////////////////////new/////////////////////////////////////////////////////////
  function new (string name, uvm_component parent);
     super.new(name, parent);
  endfunction

//////////////////////////////////////////////build_phase//////////////////////////////////////////////////////
      function void build_phase(uvm_phase phase);
		super.build_phase(phase);
   
		Rad_mon_in  = Radwa_monitor_in::type_id::create("Rad_mon_in", this);
		My_analysis_port = new("My_analysis_port", this);
	   
       $display("build phase of agent 2");
    endfunction

/////////////////////////////////////////////connect_phase/////////////////////////////////////////////////////
    function void connect_phase(uvm_phase phase);
       super.connect_phase(phase);
	   /////////////tlm
	   Rad_mon_in.analysis_port_IN.connect(My_analysis_port);
       $display("connect phase of agent 2");
    endfunction

///////////////////////////////////////////////run_phase///////////////////////////////////////////////////////
    task run_phase(uvm_phase phase);
       super.run_phase(phase);
       $display("run phase of agent 2");
    endtask

endclass

