
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////Environment/////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
class Radwa_env extends uvm_env;

  `uvm_component_utils (Radwa_env)
  
  //uvm_event monitor_done;

  Radwa_scoreboard Rad_score;
  Radwa_agent Rad_agent;
  Radwa_subscriber Rad_sub;
  Agent_IN Rad_agent_in;
  
  virtual INTF_UART U_intf;

/////////////////////////////////////////////////////new///////////////////////////////////////////////////////
  function new (string name, uvm_component parent);
  super.new(name,parent);
  endfunction
///////////////////////////////////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////build_phase/////////////////////////////////////////////////////
    function void build_phase(uvm_phase phase);
       super.build_phase(phase);
       Rad_score = Radwa_scoreboard::type_id::create("Rad_score", this);
       Rad_agent = Radwa_agent::type_id::create("Rad_agent", this);
       Rad_sub   = Radwa_subscriber::type_id::create("Rad_sub", this);
	   Rad_agent_in = Agent_IN::type_id::create("Rad_agent_in", this);

       $display("build phase of environment");
    endfunction
///////////////////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////connect_phase/////////////////////////////////////////////////////
    function void connect_phase(uvm_phase phase);
       super.connect_phase(phase);
	   ///////////////////tlm
	   /////////////////////Agent 1
	   Rad_agent.My_analysis_port.connect(Rad_sub.analysis_imp_A);
	   Rad_agent.My_analysis_port.connect(Rad_score.analysis_export_1);
	   /////////////////////Agent 2
	   Rad_agent_in.My_analysis_port.connect(Rad_sub.analysis_imp_B);
	   Rad_agent_in.My_analysis_port.connect(Rad_score.analysis_export_2);
       $display("connect phase of environment");
    endfunction
///////////////////////////////////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////run_phase////////////////////////////////////////////////////////
    task run_phase(uvm_phase phase);
       super.run_phase(phase);
       $display("run phase of environment");
    endtask
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
endclass
